** sch_path: /home/ubuntu/Desktop/design/xschem/q2_opamp_tb.sch
**.subckt q2_opamp_tb
V2 net1 net2 0 AC 0.5
V3 net1 GND 0.9
C1 OUT GND 1p m=1
.save  v(out)
V4 net3 net1 0 AC 0.5
**** begin user architecture code



.control

save all

op
write five_T_OTA_TB.raw

ac dec 10 1 10e9
set appendwrite
write five_T_OTA_TB.raw

plot db(v(out)) 180*cph(v(out))/pi

.endc



** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130B/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
**.ends
.GLOBAL GND
.end
